// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.


// Generated by Quartus Prime Version 16.0 (Build Build 211 04/27/2016)
// Created on Tue Aug 02 17:22:47 2016

module symbol_top_inst
(
//	wr_en,
	CLOCK_50,
//	data_in,
	KEY,
	VGA_HS,
	VGA_VS,
	column,
//	freeslots,
	row,
	VGA_B,
	VGA_G,
	VGA_R,
	VGA_SYNC_N,
	VGA_BLANK_N,
	VGA_CLK,
	LEDR
);

//input wire	wr_en;
input wire	CLOCK_50;
//input wire	[31:0] data_in;
input wire [3:0] KEY;
output wire	VGA_HS;
output wire	VGA_VS;
output wire	[9:0] column;
//output wire	[3:0] freeslots;
output wire	[8:0] row;
output wire	[7:0] VGA_B;
output wire	[7:0] VGA_G;
output wire	[7:0] VGA_R;
output wire [17:0] LEDR;

output wire VGA_SYNC_N, VGA_BLANK_N, VGA_CLK;

assign VGA_SYNC_N = 1'b1;
assign VGA_BLANK_N = 1'b1;

symbol_top2 u0(	// input [0:0] KEY_sig
//	.data_in(data_in) ,	// input [31:0] data_in_sig
	.KEY(KEY) ,
//	.wr_en(wr_en) ,	// input  wr_en_sig
	.CLOCK_50(CLOCK_50) ,	// input  CLOCK_50_sig
	.row(row) ,	// output [8:0] row_sig
	.column(column) ,	// output [9:0] column_sig
	.VGA_R(VGA_R) ,	// output [7:0] VGA_R_sig
	.VGA_G(VGA_G) ,	// output [7:0] VGA_G_sig
	.VGA_B(VGA_B) ,	// output [7:0] VGA_B_sig
	.VGA_HS(VGA_HS) ,	// output  VGA_HS_sig
	.VGA_VS(VGA_VS) ,	// output  VGA_VS_sig
//	.freeslots(freeslots) 	// output [3:0] freeslots_sig
	.LEDR(LEDR),
	.VGA_CLK(VGA_CLK)
	);

endmodule

