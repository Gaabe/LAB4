module resetGenerator(clkPipeline, clk, resetSig);

input clkPipeline, clk;
output resetSig;

always @(posedge clkPipeline, posedge clk)
begin
	
end

endmodule
