module S2_module(clk125, clkext, rst, sprite_number, );



endmodule
