module FIFO_writer(full, wr_en, data0, data1);

input full;
output wr_en;
output [15:0] data0, data1;

endmodule
