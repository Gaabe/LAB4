module ProcessadorGrafico()