module colisionDecoder(colisao, sp0_num, sp1_num, sp2_num, sp3_num, );

input [5:0] colisao;
input [5:0] sp0_num, sp1_num, sp2_num, sp3_num;



endmodule
