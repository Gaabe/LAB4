module mux_num2dec(sp0_num, sp1_num, sp2_num, sp3_num);



endmodule
