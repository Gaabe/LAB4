module logicLevel(logic1, logic0);

output logic1, logic0;

assign logic0 = 1'b0;
assign logic1 = 1'b1;

endmodule
